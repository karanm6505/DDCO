module demux21(input wire  a,s)